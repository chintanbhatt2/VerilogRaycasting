module FloatingPointRegister( input number [31:0]
    
);

endmodule // FloatingPointRegister